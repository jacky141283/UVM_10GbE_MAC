`ifndef TEST_LIB__SVH
`define TEST_LIB__SVH

`include "../testcases/loopback_test.sv"
`include "../testcases/packet_oversize_test.sv"

`endif
